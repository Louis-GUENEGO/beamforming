--------------------------------------------------------------------------------
--{{{ Copyright 2010 C. D. Stahl, All rights reserved.
--
--    1. Redistributions of source code must retain the above copyright 
--       notice, this list of conditions and the following disclaimer.
--    
--    2. Redistributions in binary form must reproduce the above copyright 
--       notice, this list of conditions and the following disclaimer in 
--       the documentation and/or other materials provided with the 
--       distribution.
--    
--    THIS SOFTWARE IS PROVIDED BY C. D. STAHL ``AS IS'' AND ANY EXPRESS OR 
--    IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES 
--    OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. 
--    IN NO EVENT SHALL C. D. STAHL OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, 
--    INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES 
--    (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR 
--    SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER 
--    CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT 
--    LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
--    OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF 
--    SUCH DAMAGE.
-- 
--}}}


--------------------------------------------------------------------------------
--{{{ Discription
-- This code was autogenerated by ./galois256.py.
--
-- This code describes one possible 256 element discrete field.  It includes
-- various lookup tables and functions that are common with Galois Field math.
--
-- Addition is simply xor.
--}}}


--------------------------------------------------------------------------------
--{{{ Includes
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--}}}


--------------------------------------------------------------------------------
--{{{ Package
package gf256_pkg is

  ------------------------------------------------------------------------------  
  --{{{ Types
  type gf256_map is array (natural range 0 to 255) 
    of std_logic_vector(7 downto 0);
  
  type gf256_a   is array (natural range <>) of std_logic_vector(7 downto 0);
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Zech's Logrithm
  -- This is a table mapping a power to a zech's logrithm.
  -- This can be done to perform addition in the log domain, according to the
  -- formula:
  -- a^n + a^m = a^n * (1 + a^(m-n))
  -- The zech log can be used to convert the value m-n into the value z in the
  -- below equation.
  -- a^z = (1 + a^(m-n))
  --
  -- This converts the addition into a multiplication.
  --
  --
  -- there is a special case for pwr = 00 (and pwr = FF).  In this case,
  -- (1 + a^0) = 0, which has no log representation.
  constant CONV_ZECH : gf256_map := (
    x"00", x"19", x"32", x"df", x"64", x"8a", x"bf", x"70", 
    x"c8", x"78", x"15", x"f5", x"7f", x"63", x"e0", x"21", 
    x"91", x"44", x"f0", x"5c", x"2a", x"0a", x"eb", x"c4", 
    x"fe", x"01", x"c6", x"68", x"c1", x"b5", x"42", x"2d", 
    x"23", x"0f", x"88", x"20", x"e1", x"b3", x"b8", x"6a", 
    x"54", x"9d", x"14", x"79", x"d7", x"1f", x"89", x"65", 
    x"fd", x"c5", x"02", x"ee", x"8d", x"93", x"d0", x"3f", 
    x"83", x"53", x"6b", x"52", x"84", x"ba", x"5a", x"37", 
    x"46", x"a2", x"1e", x"d8", x"11", x"82", x"40", x"6d", 
    x"c3", x"ec", x"67", x"c7", x"71", x"e4", x"d4", x"ae", 
    x"a8", x"a0", x"3b", x"39", x"28", x"aa", x"f2", x"a7", 
    x"af", x"cb", x"3e", x"d1", x"13", x"9e", x"ca", x"b0", 
    x"fb", x"be", x"8b", x"0d", x"04", x"2f", x"dd", x"4a", 
    x"1b", x"f8", x"27", x"3a", x"a1", x"47", x"7e", x"f6", 
    x"07", x"4c", x"a6", x"f3", x"d6", x"7a", x"a4", x"99", 
    x"09", x"2b", x"75", x"b7", x"b4", x"c2", x"6e", x"0c", 
    x"8c", x"ef", x"45", x"38", x"3c", x"fa", x"b1", x"90", 
    x"22", x"2e", x"05", x"62", x"80", x"34", x"da", x"96", 
    x"87", x"10", x"d9", x"35", x"ce", x"bc", x"8f", x"b2", 
    x"e2", x"77", x"c9", x"9f", x"a9", x"29", x"5d", x"9b", 
    x"51", x"6c", x"41", x"b6", x"76", x"e3", x"72", x"57", 
    x"50", x"9c", x"55", x"d3", x"e5", x"e8", x"4f", x"58", 
    x"5f", x"86", x"97", x"25", x"7c", x"1d", x"a3", x"7b", 
    x"26", x"f9", x"3d", x"cc", x"95", x"db", x"61", x"06", 
    x"f7", x"1c", x"7d", x"48", x"17", x"31", x"1a", x"4b", 
    x"08", x"9a", x"5e", x"59", x"bb", x"cf", x"94", x"cd", 
    x"36", x"5b", x"f1", x"ab", x"4e", x"e9", x"74", x"2c", 
    x"43", x"92", x"8e", x"bd", x"fc", x"66", x"ed", x"03", 
    x"0e", x"24", x"98", x"a5", x"4d", x"ac", x"e7", x"e6", 
    x"ad", x"d5", x"f4", x"16", x"49", x"de", x"33", x"81", 
    x"12", x"d2", x"56", x"73", x"ea", x"0b", x"6f", x"c0", 
    x"69", x"b9", x"85", x"60", x"dc", x"30", x"18", x"00");


  function gf256_to_zech(x : std_logic_vector)
    return std_logic_vector;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Conversion to Log
  -- This is a mapping from an element in a galois field, in polynomial form.
  -- It converts from poly to log form.  This has an issue in that there is a
  -- special case for poly = 0 mapping to a log value.  The log value is not
  -- defined for that case, but must be listed as some value.
  constant CONV_LOG : gf256_map := (
    x"00", x"00", x"01", x"19", x"02", x"32", x"1a", x"c6", 
    x"03", x"df", x"33", x"ee", x"1b", x"68", x"c7", x"4b", 
    x"04", x"64", x"e0", x"0e", x"34", x"8d", x"ef", x"81", 
    x"1c", x"c1", x"69", x"f8", x"c8", x"08", x"4c", x"71", 
    x"05", x"8a", x"65", x"2f", x"e1", x"24", x"0f", x"21", 
    x"35", x"93", x"8e", x"da", x"f0", x"12", x"82", x"45", 
    x"1d", x"b5", x"c2", x"7d", x"6a", x"27", x"f9", x"b9", 
    x"c9", x"9a", x"09", x"78", x"4d", x"e4", x"72", x"a6", 
    x"06", x"bf", x"8b", x"62", x"66", x"dd", x"30", x"fd", 
    x"e2", x"98", x"25", x"b3", x"10", x"91", x"22", x"88", 
    x"36", x"d0", x"94", x"ce", x"8f", x"96", x"db", x"bd", 
    x"f1", x"d2", x"13", x"5c", x"83", x"38", x"46", x"40", 
    x"1e", x"42", x"b6", x"a3", x"c3", x"48", x"7e", x"6e", 
    x"6b", x"3a", x"28", x"54", x"fa", x"85", x"ba", x"3d", 
    x"ca", x"5e", x"9b", x"9f", x"0a", x"15", x"79", x"2b", 
    x"4e", x"d4", x"e5", x"ac", x"73", x"f3", x"a7", x"57", 
    x"07", x"70", x"c0", x"f7", x"8c", x"80", x"63", x"0d", 
    x"67", x"4a", x"de", x"ed", x"31", x"c5", x"fe", x"18", 
    x"e3", x"a5", x"99", x"77", x"26", x"b8", x"b4", x"7c", 
    x"11", x"44", x"92", x"d9", x"23", x"20", x"89", x"2e", 
    x"37", x"3f", x"d1", x"5b", x"95", x"bc", x"cf", x"cd", 
    x"90", x"87", x"97", x"b2", x"dc", x"fc", x"be", x"61", 
    x"f2", x"56", x"d3", x"ab", x"14", x"2a", x"5d", x"9e", 
    x"84", x"3c", x"39", x"53", x"47", x"6d", x"41", x"a2", 
    x"1f", x"2d", x"43", x"d8", x"b7", x"7b", x"a4", x"76", 
    x"c4", x"17", x"49", x"ec", x"7f", x"0c", x"6f", x"f6", 
    x"6c", x"a1", x"3b", x"52", x"29", x"9d", x"55", x"aa", 
    x"fb", x"60", x"86", x"b1", x"bb", x"cc", x"3e", x"5a", 
    x"cb", x"59", x"5f", x"b0", x"9c", x"a9", x"a0", x"51", 
    x"0b", x"f5", x"16", x"eb", x"7a", x"75", x"2c", x"d7", 
    x"4f", x"ae", x"d5", x"e9", x"e6", x"e7", x"ad", x"e8", 
    x"74", x"d6", x"f4", x"ea", x"a8", x"50", x"58", x"af");


  function gf256_to_log(x : std_logic_vector)
    return std_logic_vector;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Conversion to Poly
  -- This is a mapping from the log domain to the poly domain.  There again is
  -- a special case for 0, which does not appear in this table.
  constant CONV_POLY : gf256_map := (
    x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", 
    x"1d", x"3a", x"74", x"e8", x"cd", x"87", x"13", x"26", 
    x"4c", x"98", x"2d", x"5a", x"b4", x"75", x"ea", x"c9", 
    x"8f", x"03", x"06", x"0c", x"18", x"30", x"60", x"c0", 
    x"9d", x"27", x"4e", x"9c", x"25", x"4a", x"94", x"35", 
    x"6a", x"d4", x"b5", x"77", x"ee", x"c1", x"9f", x"23", 
    x"46", x"8c", x"05", x"0a", x"14", x"28", x"50", x"a0", 
    x"5d", x"ba", x"69", x"d2", x"b9", x"6f", x"de", x"a1", 
    x"5f", x"be", x"61", x"c2", x"99", x"2f", x"5e", x"bc", 
    x"65", x"ca", x"89", x"0f", x"1e", x"3c", x"78", x"f0", 
    x"fd", x"e7", x"d3", x"bb", x"6b", x"d6", x"b1", x"7f", 
    x"fe", x"e1", x"df", x"a3", x"5b", x"b6", x"71", x"e2", 
    x"d9", x"af", x"43", x"86", x"11", x"22", x"44", x"88", 
    x"0d", x"1a", x"34", x"68", x"d0", x"bd", x"67", x"ce", 
    x"81", x"1f", x"3e", x"7c", x"f8", x"ed", x"c7", x"93", 
    x"3b", x"76", x"ec", x"c5", x"97", x"33", x"66", x"cc", 
    x"85", x"17", x"2e", x"5c", x"b8", x"6d", x"da", x"a9", 
    x"4f", x"9e", x"21", x"42", x"84", x"15", x"2a", x"54", 
    x"a8", x"4d", x"9a", x"29", x"52", x"a4", x"55", x"aa", 
    x"49", x"92", x"39", x"72", x"e4", x"d5", x"b7", x"73", 
    x"e6", x"d1", x"bf", x"63", x"c6", x"91", x"3f", x"7e", 
    x"fc", x"e5", x"d7", x"b3", x"7b", x"f6", x"f1", x"ff", 
    x"e3", x"db", x"ab", x"4b", x"96", x"31", x"62", x"c4", 
    x"95", x"37", x"6e", x"dc", x"a5", x"57", x"ae", x"41", 
    x"82", x"19", x"32", x"64", x"c8", x"8d", x"07", x"0e", 
    x"1c", x"38", x"70", x"e0", x"dd", x"a7", x"53", x"a6", 
    x"51", x"a2", x"59", x"b2", x"79", x"f2", x"f9", x"ef", 
    x"c3", x"9b", x"2b", x"56", x"ac", x"45", x"8a", x"09", 
    x"12", x"24", x"48", x"90", x"3d", x"7a", x"f4", x"f5", 
    x"f7", x"f3", x"fb", x"eb", x"cb", x"8b", x"0b", x"16", 
    x"2c", x"58", x"b0", x"7d", x"fa", x"e9", x"cf", x"83", 
    x"1b", x"36", x"6c", x"d8", x"ad", x"47", x"8e", x"01");


  function gf256_to_poly(x : std_logic_vector)
    return std_logic_vector;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Multiplicative Inverse
  -- This maps the polynomial representation of a galois field element into 
  -- another galois field element such that a^n * a^m = a^0.
  constant CONV_INV  : gf256_map := (
    x"01", x"01", x"8e", x"f4", x"47", x"a7", x"7a", x"ba", 
    x"ad", x"9d", x"dd", x"98", x"3d", x"aa", x"5d", x"96", 
    x"d8", x"72", x"c0", x"58", x"e0", x"3e", x"4c", x"66", 
    x"90", x"de", x"55", x"80", x"a0", x"83", x"4b", x"2a", 
    x"6c", x"ed", x"39", x"51", x"60", x"56", x"2c", x"8a", 
    x"70", x"d0", x"1f", x"4a", x"26", x"8b", x"33", x"6e", 
    x"48", x"89", x"6f", x"2e", x"a4", x"c3", x"40", x"5e", 
    x"50", x"22", x"cf", x"a9", x"ab", x"0c", x"15", x"e1", 
    x"36", x"5f", x"f8", x"d5", x"92", x"4e", x"a6", x"04", 
    x"30", x"88", x"2b", x"1e", x"16", x"67", x"45", x"93", 
    x"38", x"23", x"68", x"8c", x"81", x"1a", x"25", x"61", 
    x"13", x"c1", x"cb", x"63", x"97", x"0e", x"37", x"41", 
    x"24", x"57", x"ca", x"5b", x"b9", x"c4", x"17", x"4d", 
    x"52", x"8d", x"ef", x"b3", x"20", x"ec", x"2f", x"32", 
    x"28", x"d1", x"11", x"d9", x"e9", x"fb", x"da", x"79", 
    x"db", x"77", x"06", x"bb", x"84", x"cd", x"fe", x"fc", 
    x"1b", x"54", x"a1", x"1d", x"7c", x"cc", x"e4", x"b0", 
    x"49", x"31", x"27", x"2d", x"53", x"69", x"02", x"f5", 
    x"18", x"df", x"44", x"4f", x"9b", x"bc", x"0f", x"5c", 
    x"0b", x"dc", x"bd", x"94", x"ac", x"09", x"c7", x"a2", 
    x"1c", x"82", x"9f", x"c6", x"34", x"c2", x"46", x"05", 
    x"ce", x"3b", x"0d", x"3c", x"9c", x"08", x"be", x"b7", 
    x"87", x"e5", x"ee", x"6b", x"eb", x"f2", x"bf", x"af", 
    x"c5", x"64", x"07", x"7b", x"95", x"9a", x"ae", x"b6", 
    x"12", x"59", x"a5", x"35", x"65", x"b8", x"a3", x"9e", 
    x"d2", x"f7", x"62", x"5a", x"85", x"7d", x"a8", x"3a", 
    x"29", x"71", x"c8", x"f6", x"f9", x"43", x"d7", x"d6", 
    x"10", x"73", x"76", x"78", x"99", x"0a", x"19", x"91", 
    x"14", x"3f", x"e6", x"f0", x"86", x"b1", x"e2", x"f1", 
    x"fa", x"74", x"f3", x"b4", x"6d", x"21", x"b2", x"6a", 
    x"e3", x"e7", x"b5", x"ea", x"03", x"8f", x"d3", x"c9", 
    x"42", x"d4", x"e8", x"75", x"7f", x"ff", x"7e", x"fd");


  function gf256_invert(x : std_logic_vector)
    return std_logic_vector;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Galois Field Multiply
  function gf256_mult(x : std_logic_vector; y : std_logic_vector)
    return std_logic_vector;
  --}}}


end package;
--}}}


-------------------------------------------------------------------------------
--{{{ Package Body
package body gf256_pkg is

  ------------------------------------------------------------------------------
  --{{{ Zech's Logrithm
  function gf256_to_zech(x : std_logic_vector)
      return std_logic_vector is
  begin
    return CONV_ZECH(to_integer(unsigned(x)));
  end function;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Conversion to Log
  function gf256_to_log(x : std_logic_vector)
      return std_logic_vector is
  begin
    return CONV_LOG(to_integer(unsigned(x)));
  end function;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Conversion to Poly
  function gf256_to_poly(x : std_logic_vector)
      return std_logic_vector is
  begin
    return CONV_POLY(to_integer(unsigned(x)));
  end function;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Multiplicative Inverse
  function gf256_invert(x : std_logic_vector)
      return std_logic_vector is
  begin
    return CONV_INV(to_integer(unsigned(x)));
  end function;
  --}}}


  ------------------------------------------------------------------------------
  --{{{ Galois Field Multiply
  function gf256_mult(x : std_logic_vector; y : std_logic_vector)
      return std_logic_vector is
    variable tmp : std_logic_vector(7 downto 0);
  begin
    tmp(0) := (x(6) and y(2)) xor (x(3) and y(5)) xor (x(4) and y(4))
              xor (x(5) and y(3)) xor (x(0) and y(0)) xor (x(5) and y(7))
              xor (x(7) and y(6)) xor (x(7) and y(7)) xor (x(1) and y(7))
              xor (x(7) and y(5)) xor (x(7) and y(1)) xor (x(2) and y(6))
              xor (x(6) and y(7)) xor (x(6) and y(6));
    tmp(1) := (x(3) and y(6)) xor (x(0) and y(1)) xor (x(4) and y(5))
              xor (x(7) and y(6)) xor (x(7) and y(2)) xor (x(5) and y(4))
              xor (x(7) and y(7)) xor (x(1) and y(0)) xor (x(6) and y(3))
              xor (x(2) and y(7)) xor (x(6) and y(7));
    tmp(2) := (x(6) and y(4)) xor (x(7) and y(3)) xor (x(4) and y(6))
              xor (x(4) and y(4)) xor (x(5) and y(3)) xor (x(3) and y(7))
              xor (x(5) and y(7)) xor (x(7) and y(6)) xor (x(1) and y(1))
              xor (x(1) and y(7)) xor (x(7) and y(5)) xor (x(3) and y(5))
              xor (x(7) and y(1)) xor (x(2) and y(6)) xor (x(5) and y(5))
              xor (x(6) and y(2)) xor (x(6) and y(6)) xor (x(2) and y(0))
              xor (x(6) and y(7)) xor (x(0) and y(2));
    tmp(3) := (x(0) and y(3)) xor (x(7) and y(4)) xor (x(1) and y(2))
              xor (x(7) and y(5)) xor (x(5) and y(4)) xor (x(2) and y(1))
              xor (x(2) and y(7)) xor (x(2) and y(6)) xor (x(6) and y(5))
              xor (x(6) and y(3)) xor (x(6) and y(6)) xor (x(6) and y(2))
              xor (x(4) and y(7)) xor (x(4) and y(5)) xor (x(4) and y(4))
              xor (x(7) and y(1)) xor (x(3) and y(6)) xor (x(5) and y(6))
              xor (x(5) and y(7)) xor (x(1) and y(7)) xor (x(3) and y(0))
              xor (x(3) and y(5)) xor (x(5) and y(3)) xor (x(7) and y(2));
    tmp(4) := (x(0) and y(4)) xor (x(7) and y(7)) xor (x(1) and y(7))
              xor (x(7) and y(3)) xor (x(3) and y(1)) xor (x(2) and y(7))
              xor (x(2) and y(6)) xor (x(6) and y(4)) xor (x(4) and y(0))
              xor (x(4) and y(6)) xor (x(4) and y(5)) xor (x(4) and y(4))
              xor (x(5) and y(3)) xor (x(7) and y(2)) xor (x(3) and y(7))
              xor (x(5) and y(4)) xor (x(5) and y(5)) xor (x(2) and y(2))
              xor (x(6) and y(3)) xor (x(1) and y(3)) xor (x(6) and y(2))
              xor (x(3) and y(5)) xor (x(7) and y(1)) xor (x(3) and y(6));
    tmp(5) := (x(3) and y(6)) xor (x(0) and y(5)) xor (x(7) and y(3))
              xor (x(7) and y(4)) xor (x(1) and y(4)) xor (x(3) and y(2))
              xor (x(6) and y(3)) xor (x(5) and y(4)) xor (x(6) and y(5))
              xor (x(6) and y(4)) xor (x(4) and y(1)) xor (x(4) and y(7))
              xor (x(4) and y(6)) xor (x(4) and y(5)) xor (x(5) and y(0))
              xor (x(3) and y(7)) xor (x(5) and y(6)) xor (x(2) and y(3))
              xor (x(5) and y(5)) xor (x(2) and y(7)) xor (x(7) and y(2));
    tmp(6) := (x(4) and y(2)) xor (x(3) and y(7)) xor (x(5) and y(1))
              xor (x(4) and y(7)) xor (x(4) and y(6)) xor (x(0) and y(6))
              xor (x(7) and y(5)) xor (x(5) and y(6)) xor (x(1) and y(5))
              xor (x(7) and y(4)) xor (x(5) and y(7)) xor (x(3) and y(3))
              xor (x(2) and y(4)) xor (x(6) and y(0)) xor (x(5) and y(5))
              xor (x(6) and y(5)) xor (x(6) and y(4)) xor (x(7) and y(3))
              xor (x(6) and y(6));
    tmp(7) := (x(4) and y(3)) xor (x(5) and y(2)) xor (x(4) and y(7))
              xor (x(3) and y(4)) xor (x(7) and y(0)) xor (x(5) and y(6))
              xor (x(7) and y(4)) xor (x(5) and y(7)) xor (x(0) and y(7))
              xor (x(7) and y(5)) xor (x(2) and y(5)) xor (x(7) and y(6))
              xor (x(1) and y(6)) xor (x(6) and y(1)) xor (x(6) and y(5))
              xor (x(6) and y(7)) xor (x(6) and y(6));

    return tmp;
  end function;
  --}}}

end package body;
--}}}

